library IEEE; 
use IEEE.STD_LOGIC_1164.all; 

package mypackage is 

   
        type ops is (ADD, SUB, ZERO, SHR, SHL, NOP, ROL_O, ROR_O, INC, DEC);

end mypackage; 


